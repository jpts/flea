magic
tech scmos
timestamp 695379524
<< polysilicon >>
rect -26 -2 25 4
<< metal1 >>
rect 20 -3 25 5
<< labels >>
rlabel metal1 23 1 23 1 7 right
rlabel polysilicon -24 1 -24 1 3 left
rlabel space -2 10 -2 10 5 top
rlabel space -1 -5 -1 -5 1 bottom
<< end >>
