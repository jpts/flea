magic
tech scmos
timestamp 597519242
<< polysilicon >>
rect -24 269 -22 270
rect -24 267 -19 269
rect 173 267 175 269
rect 101 238 121 240
rect 101 235 105 238
rect 130 235 138 237
rect -6 210 -4 214
rect 10 210 13 214
rect 17 210 27 214
rect 41 210 43 214
rect -6 192 -4 196
rect 10 193 13 196
rect 17 193 27 196
rect 10 192 27 193
rect 41 192 43 196
rect 19 189 25 192
rect -6 160 -4 164
rect 10 160 20 164
rect 24 160 27 164
rect 41 160 43 164
rect -6 142 -4 146
rect 10 142 20 146
rect 24 142 27 146
rect 41 142 43 146
rect 12 139 18 142
rect -17 125 -15 128
rect 101 219 105 221
rect 130 219 138 221
rect 82 201 86 203
rect 132 201 136 219
rect 341 212 343 215
rect 170 210 343 212
rect 170 208 172 210
rect 170 206 343 208
rect 82 190 86 194
rect 132 190 136 194
rect 82 173 86 183
rect 100 173 104 175
rect 132 173 136 183
rect 150 173 154 175
rect 82 156 86 166
rect 100 164 104 166
rect 100 158 107 164
rect 132 163 136 166
rect 100 156 104 158
rect 103 152 104 156
rect 82 149 86 152
rect 100 149 104 152
rect 132 149 136 159
rect 150 163 154 166
rect 150 149 154 159
rect 82 140 86 142
rect 100 140 104 142
rect 132 140 136 142
rect 150 140 154 142
rect 341 204 343 206
rect 170 202 343 204
rect 170 200 172 202
rect 170 198 343 200
rect 341 196 343 198
rect 170 194 343 196
rect 170 192 172 194
rect 170 190 343 192
rect 341 188 343 190
rect 170 186 343 188
rect 170 184 172 186
rect 170 182 343 184
rect 341 180 343 182
rect 170 178 343 180
rect 170 176 172 178
rect 170 174 343 176
rect 341 172 343 174
rect 170 170 343 172
rect 170 168 172 170
rect 170 166 343 168
rect 341 164 343 166
rect 170 162 343 164
rect 170 160 172 162
rect 170 158 343 160
rect 341 156 343 158
rect 170 154 343 156
rect 170 152 172 154
rect 170 150 343 152
rect 341 148 343 150
rect 170 146 343 148
rect 170 144 172 146
rect 170 142 343 144
rect 341 140 343 142
rect 170 138 343 140
rect 170 136 172 138
rect 170 134 343 136
rect 341 132 343 134
rect 170 130 343 132
rect 170 128 172 130
rect 170 126 343 128
rect -17 123 156 125
rect 154 121 156 123
rect 341 124 343 126
rect 166 122 343 124
rect -17 119 156 121
rect -17 116 -15 119
<< ndiffusion >>
rect 100 221 101 235
rect 105 221 106 235
rect 129 221 130 235
rect 138 221 139 235
rect 81 194 82 201
rect 86 194 87 201
rect 131 194 132 201
rect 136 194 137 201
rect 81 183 82 190
rect 86 183 87 190
rect 131 183 132 190
rect 136 183 137 190
rect 81 166 82 173
rect 86 166 87 173
rect 99 166 100 173
rect 104 166 105 173
rect 131 166 132 173
rect 136 166 137 173
rect 149 166 150 173
rect 154 166 155 173
rect 81 142 82 149
rect 86 142 87 149
rect 99 142 100 149
rect 104 142 105 149
rect 131 142 132 149
rect 136 142 137 149
rect 149 142 150 149
rect 154 142 155 149
rect 15 99 33 103
rect 15 95 19 99
rect 23 95 33 99
rect 15 91 33 95
rect 59 99 77 103
rect 59 95 63 99
rect 67 95 77 99
rect 59 91 77 95
rect 103 99 121 103
rect 103 95 107 99
rect 111 95 121 99
rect 103 91 121 95
rect 147 99 165 103
rect 147 95 151 99
rect 155 95 165 99
rect 147 91 165 95
rect 191 99 209 103
rect 191 95 195 99
rect 199 95 209 99
rect 191 91 209 95
rect 15 61 33 65
rect 15 57 19 61
rect 23 57 33 61
rect 15 53 33 57
rect 59 61 77 65
rect 59 57 63 61
rect 67 57 77 61
rect 59 53 77 57
rect 103 61 121 65
rect 103 57 107 61
rect 111 57 121 61
rect 103 53 121 57
rect 147 61 165 65
rect 147 57 151 61
rect 155 57 165 61
rect 147 53 165 57
rect 191 61 209 65
rect 191 57 195 61
rect 199 57 209 61
rect 191 53 209 57
rect 235 61 253 65
rect 235 57 239 61
rect 243 57 253 61
rect 235 53 253 57
rect 15 23 33 27
rect 15 19 19 23
rect 23 19 33 23
rect 15 15 33 19
rect 59 23 77 27
rect 59 19 63 23
rect 67 19 77 23
rect 59 15 77 19
rect 103 23 121 27
rect 103 19 107 23
rect 111 19 121 23
rect 103 15 121 19
rect 147 23 165 27
rect 147 19 151 23
rect 155 19 165 23
rect 147 15 165 19
rect 191 23 209 27
rect 191 19 195 23
rect 199 19 209 23
rect 191 15 209 19
rect 235 23 253 27
rect 235 19 239 23
rect 243 19 253 23
rect 235 15 253 19
<< pdiffusion >>
rect -19 269 173 270
rect -19 266 173 267
rect -4 214 10 215
rect 27 214 41 215
rect -4 209 10 210
rect 27 209 41 210
rect -4 196 10 197
rect 27 196 41 197
rect -4 191 10 192
rect 27 191 41 192
rect -4 164 10 165
rect 27 164 41 165
rect -4 159 10 160
rect 27 159 41 160
rect -4 146 10 147
rect 27 146 41 147
rect -4 141 10 142
rect 27 141 41 142
<< metal1 >>
rect -26 274 -22 280
rect 178 279 182 280
rect -22 270 -19 274
rect -26 256 -22 270
rect -26 252 -19 256
rect -29 136 -19 140
rect -15 252 -13 256
rect 71 241 75 242
rect 13 233 68 236
rect 13 224 17 233
rect 5 219 9 220
rect 13 214 17 220
rect -11 205 -4 209
rect -11 201 -7 205
rect 13 201 17 210
rect 10 197 17 201
rect 20 227 62 230
rect 20 209 24 227
rect 27 219 31 220
rect 41 205 48 209
rect 20 201 24 205
rect 20 197 27 201
rect -11 181 -7 197
rect 24 190 27 191
rect 10 187 11 190
rect 20 187 27 190
rect 44 186 48 205
rect 44 181 48 182
rect -11 178 17 181
rect 6 169 10 170
rect 13 159 17 178
rect -11 155 -4 159
rect -11 136 -7 155
rect 13 151 17 155
rect 10 147 17 151
rect 20 178 48 181
rect 20 174 24 178
rect 20 164 24 170
rect 28 169 32 170
rect 20 151 24 160
rect 41 155 48 159
rect 44 151 48 155
rect 20 147 27 151
rect 20 146 24 147
rect 10 140 13 141
rect 10 137 17 140
rect -29 90 -25 136
rect 27 136 31 137
rect 44 128 48 147
rect -18 125 48 128
rect 59 156 62 227
rect 65 224 68 233
rect 106 235 110 242
rect 65 221 96 224
rect 125 235 129 262
rect 178 256 182 257
rect 182 252 351 256
rect 163 241 167 242
rect 110 221 111 225
rect 143 221 151 225
rect 155 221 163 225
rect 167 222 351 226
rect 167 221 171 222
rect 65 163 68 221
rect 78 215 340 218
rect 344 215 351 219
rect 78 201 81 215
rect 131 206 137 210
rect 137 201 141 206
rect 77 190 81 194
rect 87 190 131 194
rect 137 190 141 194
rect 137 180 141 183
rect 163 205 167 206
rect 87 176 110 180
rect 114 176 118 180
rect 87 173 91 176
rect 76 166 77 170
rect 95 163 99 166
rect 105 163 109 166
rect 65 159 87 163
rect 91 159 99 163
rect 106 159 109 163
rect 115 163 118 176
rect 137 176 163 180
rect 137 173 141 176
rect 155 173 163 176
rect 126 167 127 171
rect 159 166 163 173
rect 145 163 149 166
rect 115 159 122 163
rect 126 159 132 163
rect 136 159 150 163
rect 59 152 72 156
rect 76 152 82 156
rect 86 152 99 156
rect 95 149 99 152
rect 115 152 137 156
rect 141 152 149 156
rect 106 149 109 150
rect 76 144 77 148
rect 87 139 91 142
rect 115 139 118 152
rect 145 149 149 152
rect 157 149 163 166
rect 126 145 127 149
rect 159 142 163 149
rect 87 135 95 139
rect 99 135 118 139
rect 137 139 141 142
rect 155 139 163 142
rect 137 133 163 139
rect 137 132 167 133
rect 52 118 56 127
rect 161 121 162 125
rect -18 99 -14 112
rect 0 113 4 114
rect -29 86 0 90
rect 44 113 48 114
rect 4 104 10 108
rect 38 104 44 108
rect 4 103 14 104
rect 4 91 10 103
rect 34 103 44 104
rect 23 95 25 99
rect 4 90 14 91
rect 38 91 44 103
rect 34 90 44 91
rect 4 86 10 90
rect 38 86 44 90
rect 0 80 4 81
rect 88 113 92 114
rect 48 104 54 108
rect 82 104 88 108
rect 48 103 58 104
rect 48 91 54 103
rect 78 103 88 104
rect 67 95 69 99
rect 48 90 58 91
rect 82 91 88 103
rect 78 90 88 91
rect 48 86 54 90
rect 82 86 88 90
rect 44 80 48 81
rect 132 113 136 114
rect 92 104 98 108
rect 126 104 132 108
rect 92 103 102 104
rect 92 91 98 103
rect 122 103 132 104
rect 111 95 113 99
rect 92 90 102 91
rect 126 91 132 103
rect 122 90 132 91
rect 92 86 98 90
rect 126 86 132 90
rect 88 80 92 81
rect 176 113 180 114
rect 136 104 142 108
rect 170 104 176 108
rect 136 103 146 104
rect 136 91 142 103
rect 166 103 176 104
rect 155 95 157 99
rect 136 90 146 91
rect 170 91 176 103
rect 166 90 176 91
rect 136 86 142 90
rect 170 86 176 90
rect 132 80 136 81
rect 220 113 224 114
rect 180 104 186 108
rect 214 104 220 108
rect 180 103 190 104
rect 180 91 186 103
rect 210 103 220 104
rect 199 95 201 99
rect 180 90 190 91
rect 214 91 220 103
rect 210 90 220 91
rect 180 86 186 90
rect 214 86 220 90
rect 176 80 180 81
rect 220 80 224 81
rect 0 75 4 76
rect 44 75 48 76
rect 4 66 10 70
rect 38 66 44 70
rect 4 65 14 66
rect 4 53 10 65
rect 34 65 44 66
rect 23 57 25 61
rect 4 52 14 53
rect 38 53 44 65
rect 34 52 44 53
rect 4 48 10 52
rect 38 48 44 52
rect 0 42 4 43
rect 88 75 92 76
rect 48 66 54 70
rect 82 66 88 70
rect 48 65 58 66
rect 48 53 54 65
rect 78 65 88 66
rect 67 57 69 61
rect 48 52 58 53
rect 82 53 88 65
rect 78 52 88 53
rect 48 48 54 52
rect 82 48 88 52
rect 44 42 48 43
rect 132 75 136 76
rect 92 66 98 70
rect 126 66 132 70
rect 92 65 102 66
rect 92 53 98 65
rect 122 65 132 66
rect 111 57 113 61
rect 92 52 102 53
rect 126 53 132 65
rect 122 52 132 53
rect 92 48 98 52
rect 126 48 132 52
rect 88 42 92 43
rect 176 75 180 76
rect 136 66 142 70
rect 170 66 176 70
rect 136 65 146 66
rect 136 53 142 65
rect 166 65 176 66
rect 155 57 157 61
rect 136 52 146 53
rect 170 53 176 65
rect 166 52 176 53
rect 136 48 142 52
rect 170 48 176 52
rect 132 42 136 43
rect 220 75 224 76
rect 180 66 186 70
rect 214 66 220 70
rect 180 65 190 66
rect 180 53 186 65
rect 210 65 220 66
rect 199 57 201 61
rect 180 52 190 53
rect 214 53 220 65
rect 210 52 220 53
rect 180 48 186 52
rect 214 48 220 52
rect 176 42 180 43
rect 264 75 268 76
rect 224 66 230 70
rect 258 66 264 70
rect 224 65 234 66
rect 224 53 230 65
rect 254 65 264 66
rect 243 57 245 61
rect 224 52 234 53
rect 258 53 264 65
rect 254 52 264 53
rect 224 48 230 52
rect 258 48 264 52
rect 220 42 224 43
rect 264 42 268 43
rect 0 37 4 38
rect 44 37 48 38
rect 4 28 10 32
rect 38 28 44 32
rect 4 27 14 28
rect 4 15 10 27
rect 34 27 44 28
rect 23 19 25 23
rect 4 14 14 15
rect 38 15 44 27
rect 34 14 44 15
rect 4 10 10 14
rect 38 10 44 14
rect 0 4 4 5
rect 88 37 92 38
rect 48 28 54 32
rect 82 28 88 32
rect 48 27 58 28
rect 48 15 54 27
rect 78 27 88 28
rect 67 19 69 23
rect 48 14 58 15
rect 82 15 88 27
rect 78 14 88 15
rect 48 10 54 14
rect 82 10 88 14
rect 44 4 48 5
rect 132 37 136 38
rect 92 28 98 32
rect 126 28 132 32
rect 92 27 102 28
rect 92 15 98 27
rect 122 27 132 28
rect 111 19 113 23
rect 92 14 102 15
rect 126 15 132 27
rect 122 14 132 15
rect 92 10 98 14
rect 126 10 132 14
rect 88 4 92 5
rect 176 37 180 38
rect 136 28 142 32
rect 170 28 176 32
rect 136 27 146 28
rect 136 15 142 27
rect 166 27 176 28
rect 155 19 157 23
rect 136 14 146 15
rect 170 15 176 27
rect 166 14 176 15
rect 136 10 142 14
rect 170 10 176 14
rect 132 4 136 5
rect 220 37 224 38
rect 180 28 186 32
rect 214 28 220 32
rect 180 27 190 28
rect 180 15 186 27
rect 210 27 220 28
rect 199 19 201 23
rect 180 14 190 15
rect 214 15 220 27
rect 210 14 220 15
rect 180 10 186 14
rect 214 10 220 14
rect 176 4 180 5
rect 264 37 268 38
rect 224 28 230 32
rect 258 28 264 32
rect 224 27 234 28
rect 224 15 230 27
rect 254 27 264 28
rect 243 19 245 23
rect 224 14 234 15
rect 258 15 264 27
rect 254 14 264 15
rect 224 10 230 14
rect 258 10 264 14
rect 220 4 224 5
rect 264 4 268 5
<< metal2 >>
rect 17 220 27 224
rect 5 209 9 220
rect 111 210 115 221
rect 5 205 20 209
rect 151 210 155 221
rect -7 197 24 201
rect 20 194 24 197
rect 11 182 44 186
rect 110 180 352 181
rect 114 176 352 180
rect 10 170 20 174
rect 28 159 32 170
rect 17 155 32 159
rect 72 156 76 166
rect 13 147 44 151
rect 87 148 91 159
rect 13 144 17 147
rect 76 144 91 148
rect 95 159 102 163
rect 95 139 99 159
rect 110 150 114 176
rect 126 167 141 171
rect 122 149 126 159
rect 137 156 141 167
rect -7 132 27 136
rect 31 132 48 136
rect -14 95 25 99
rect 25 61 29 95
rect 44 61 48 132
rect 157 99 161 121
rect 73 95 113 99
rect 113 61 117 95
rect 44 57 69 61
rect 25 23 29 57
rect 113 23 117 57
rect 29 19 69 23
rect 73 19 113 23
rect 157 61 161 95
rect 201 61 205 95
rect 205 57 245 61
rect 157 23 161 57
rect 245 23 249 57
rect 161 19 201 23
rect 205 19 245 23
<< pwell >>
rect 71 210 167 246
rect 65 128 167 210
rect 10 86 38 108
rect 54 86 82 108
rect 98 86 126 108
rect 142 86 170 108
rect 186 86 214 108
rect 10 48 38 70
rect 54 48 82 70
rect 98 48 126 70
rect 142 48 170 70
rect 186 48 214 70
rect 230 48 258 70
rect 10 10 38 32
rect 54 10 82 32
rect 98 10 126 32
rect 142 10 170 32
rect 186 10 214 32
rect 230 10 258 32
<< polycontact >>
rect -26 270 -22 274
rect 121 237 125 241
rect 13 210 17 214
rect 13 193 17 197
rect 20 160 24 164
rect 20 142 24 146
rect -18 128 -14 132
rect 340 215 344 219
rect 132 159 136 163
rect 82 152 86 156
rect 99 152 103 156
rect 150 159 154 163
rect 162 121 166 125
rect -18 112 -14 116
<< ndcontact >>
rect 96 221 100 235
rect 106 221 110 235
rect 125 221 129 235
rect 139 221 143 235
rect 77 194 81 201
rect 87 194 91 201
rect 127 194 131 201
rect 137 194 141 201
rect 77 183 81 190
rect 87 183 91 190
rect 127 183 131 190
rect 137 183 141 190
rect 77 166 81 173
rect 87 166 91 173
rect 95 166 99 173
rect 105 166 109 173
rect 127 166 131 173
rect 137 166 141 173
rect 145 166 149 173
rect 155 166 159 173
rect 77 142 81 149
rect 87 142 91 149
rect 95 142 99 149
rect 105 142 109 149
rect 127 142 131 149
rect 137 142 141 149
rect 145 142 149 149
rect 155 142 159 149
rect 19 95 23 99
rect 63 95 67 99
rect 107 95 111 99
rect 151 95 155 99
rect 195 95 199 99
rect 19 57 23 61
rect 63 57 67 61
rect 107 57 111 61
rect 151 57 155 61
rect 195 57 199 61
rect 239 57 243 61
rect 19 19 23 23
rect 63 19 67 23
rect 107 19 111 23
rect 151 19 155 23
rect 195 19 199 23
rect 239 19 243 23
<< pdcontact >>
rect -19 270 173 274
rect -19 262 173 266
rect -4 215 10 219
rect 27 215 41 219
rect -4 205 10 209
rect 27 205 41 209
rect -4 197 10 201
rect 27 197 41 201
rect -4 187 10 191
rect 27 187 41 191
rect -4 165 10 169
rect 27 165 41 169
rect -4 155 10 159
rect 27 155 41 159
rect -4 147 10 151
rect 27 147 41 151
rect -4 137 10 141
rect 27 137 41 141
<< m2contact >>
rect 5 220 9 224
rect 13 220 17 224
rect -11 197 -7 201
rect 27 220 31 224
rect 20 205 24 209
rect 20 190 24 194
rect 11 186 15 190
rect 44 182 48 186
rect 6 170 10 174
rect 13 155 17 159
rect 20 170 24 174
rect 28 170 32 174
rect 44 147 48 151
rect 13 140 17 144
rect -11 132 -7 136
rect 27 132 31 136
rect 111 221 115 225
rect 151 221 155 225
rect 111 206 115 210
rect 151 206 155 210
rect 110 176 114 180
rect 72 166 76 170
rect 87 159 91 163
rect 102 159 106 163
rect 122 167 126 171
rect 122 159 126 163
rect 72 152 76 156
rect 106 150 110 154
rect 137 152 141 156
rect 72 144 76 148
rect 122 145 126 149
rect 95 135 99 139
rect 157 121 161 125
rect -18 95 -14 99
rect 25 95 29 99
rect 69 95 73 99
rect 113 95 117 99
rect 157 95 161 99
rect 201 95 205 99
rect 25 57 29 61
rect 69 57 73 61
rect 113 57 117 61
rect 157 57 161 61
rect 201 57 205 61
rect 245 57 249 61
rect 25 19 29 23
rect 69 19 73 23
rect 113 19 117 23
rect 157 19 161 23
rect 201 19 205 23
rect 245 19 249 23
<< ntransistor >>
rect 101 221 105 235
rect 130 221 138 235
rect 82 194 86 201
rect 132 194 136 201
rect 82 183 86 190
rect 132 183 136 190
rect 82 166 86 173
rect 100 166 104 173
rect 132 166 136 173
rect 150 166 154 173
rect 82 142 86 149
rect 100 142 104 149
rect 132 142 136 149
rect 150 142 154 149
<< ptransistor >>
rect -19 267 173 269
rect -4 210 10 214
rect 27 210 41 214
rect -4 192 10 196
rect 27 192 41 196
rect -4 160 10 164
rect 27 160 41 164
rect -4 142 10 146
rect 27 142 41 146
<< psubstratepcontact >>
rect 71 242 118 246
rect 133 242 167 246
rect 71 227 75 241
rect 163 221 167 241
rect 84 206 111 210
rect 115 206 131 210
rect 137 206 151 210
rect 155 206 167 210
rect 163 133 167 205
rect 68 128 167 132
rect 10 104 38 108
rect 10 91 14 103
rect 34 91 38 103
rect 10 86 38 90
rect 54 104 82 108
rect 54 91 58 103
rect 78 91 82 103
rect 54 86 82 90
rect 98 104 126 108
rect 98 91 102 103
rect 122 91 126 103
rect 98 86 126 90
rect 142 104 170 108
rect 142 91 146 103
rect 166 91 170 103
rect 142 86 170 90
rect 186 104 214 108
rect 186 91 190 103
rect 210 91 214 103
rect 186 86 214 90
rect 10 66 38 70
rect 10 53 14 65
rect 34 53 38 65
rect 10 48 38 52
rect 54 66 82 70
rect 54 53 58 65
rect 78 53 82 65
rect 54 48 82 52
rect 98 66 126 70
rect 98 53 102 65
rect 122 53 126 65
rect 98 48 126 52
rect 142 66 170 70
rect 142 53 146 65
rect 166 53 170 65
rect 142 48 170 52
rect 186 66 214 70
rect 186 53 190 65
rect 210 53 214 65
rect 186 48 214 52
rect 230 66 258 70
rect 230 53 234 65
rect 254 53 258 65
rect 230 48 258 52
rect 10 28 38 32
rect 10 15 14 27
rect 34 15 38 27
rect 10 10 38 14
rect 54 28 82 32
rect 54 15 58 27
rect 78 15 82 27
rect 54 10 82 14
rect 98 28 126 32
rect 98 15 102 27
rect 122 15 126 27
rect 98 10 126 14
rect 142 28 170 32
rect 142 15 146 27
rect 166 15 170 27
rect 142 10 170 14
rect 186 28 214 32
rect 186 15 190 27
rect 210 15 214 27
rect 186 10 214 14
rect 230 28 258 32
rect 230 15 234 27
rect 254 15 258 27
rect 230 10 258 14
<< nsubstratencontact >>
rect -26 280 182 284
rect 178 257 182 279
rect -19 136 -15 256
rect -13 252 121 256
rect 133 252 182 256
rect 52 127 56 222
rect 0 114 224 118
rect 0 81 4 113
rect 44 81 48 113
rect 88 81 92 113
rect 132 81 136 113
rect 176 81 180 113
rect 220 81 224 113
rect 0 76 268 80
rect 0 43 4 75
rect 44 43 48 75
rect 88 43 92 75
rect 132 43 136 75
rect 176 43 180 75
rect 220 43 224 75
rect 264 43 268 75
rect 0 38 268 42
rect 0 5 4 37
rect 44 5 48 37
rect 88 5 92 37
rect 132 5 136 37
rect 176 5 180 37
rect 220 5 224 37
rect 264 5 268 37
rect 0 0 268 4
<< psubstratepdiff >>
rect 118 242 133 246
rect 71 241 75 242
rect 163 241 167 242
rect 71 210 75 227
rect 110 210 116 211
rect 65 206 84 210
rect 111 206 115 210
rect 65 132 69 206
rect 110 205 116 206
rect 150 210 156 211
rect 163 210 167 221
rect 151 206 155 210
rect 150 205 156 206
rect 163 205 167 206
rect 163 132 167 133
rect 65 128 68 132
rect 10 103 38 104
rect 14 91 15 103
rect 33 91 34 103
rect 10 90 38 91
rect 54 103 82 104
rect 58 91 59 103
rect 77 91 78 103
rect 54 90 82 91
rect 98 103 126 104
rect 102 91 103 103
rect 121 91 122 103
rect 98 90 126 91
rect 142 103 170 104
rect 146 91 147 103
rect 165 91 166 103
rect 142 90 170 91
rect 186 103 214 104
rect 190 91 191 103
rect 209 91 210 103
rect 186 90 214 91
rect 10 65 38 66
rect 14 53 15 65
rect 33 53 34 65
rect 10 52 38 53
rect 54 65 82 66
rect 58 53 59 65
rect 77 53 78 65
rect 54 52 82 53
rect 98 65 126 66
rect 102 53 103 65
rect 121 53 122 65
rect 98 52 126 53
rect 142 65 170 66
rect 146 53 147 65
rect 165 53 166 65
rect 142 52 170 53
rect 186 65 214 66
rect 190 53 191 65
rect 209 53 210 65
rect 186 52 214 53
rect 230 65 258 66
rect 234 53 235 65
rect 253 53 254 65
rect 230 52 258 53
rect 10 27 38 28
rect 14 15 15 27
rect 33 15 34 27
rect 10 14 38 15
rect 54 27 82 28
rect 58 15 59 27
rect 77 15 78 27
rect 54 14 82 15
rect 98 27 126 28
rect 102 15 103 27
rect 121 15 122 27
rect 98 14 126 15
rect 142 27 170 28
rect 146 15 147 27
rect 165 15 166 27
rect 142 14 170 15
rect 186 27 214 28
rect 190 15 191 27
rect 209 15 210 27
rect 186 14 214 15
rect 230 27 258 28
rect 234 15 235 27
rect 253 15 254 27
rect 230 14 258 15
<< nsubstratendiff >>
rect 178 279 182 280
rect 178 256 182 257
rect -15 252 -13 256
rect 0 113 4 114
rect 44 113 48 114
rect 0 80 4 81
rect 88 113 92 114
rect 44 80 48 81
rect 132 113 136 114
rect 88 80 92 81
rect 176 113 180 114
rect 132 80 136 81
rect 220 113 224 114
rect 176 80 180 81
rect 220 80 224 81
rect 0 75 4 76
rect 44 75 48 76
rect 0 42 4 43
rect 88 75 92 76
rect 44 42 48 43
rect 132 75 136 76
rect 88 42 92 43
rect 176 75 180 76
rect 132 42 136 43
rect 220 75 224 76
rect 176 42 180 43
rect 264 75 268 76
rect 220 42 224 43
rect 264 42 268 43
rect 0 37 4 38
rect 44 37 48 38
rect 0 4 4 5
rect 88 37 92 38
rect 44 4 48 5
rect 132 37 136 38
rect 88 4 92 5
rect 176 37 180 38
rect 132 4 136 5
rect 220 37 224 38
rect 176 4 180 5
rect 264 37 268 38
rect 220 4 224 5
rect 264 4 268 5
<< labels >>
rlabel ptransistor -4 160 10 164 0 m1
rlabel ptransistor 27 142 41 146 0 m1
rlabel ptransistor 27 160 41 164 0 m2
rlabel ptransistor -4 142 10 146 0 m2
rlabel metal1 46 129 46 129 1 node10
rlabel metal1 15 177 15 177 1 node7
rlabel metal1 22 177 22 177 1 node8
rlabel ptransistor 27 210 41 214 0 m3
rlabel ptransistor -4 192 10 196 0 m3
rlabel ptransistor -4 210 10 214 0 m4
rlabel ptransistor 27 192 41 196 0 m4
rlabel metal1 79 213 79 213 1 node13
rlabel pwell 112 192 112 192 1 node14
rlabel ntransistor 82 194 86 201 0 m10
rlabel ntransistor 82 183 86 190 0 m10
rlabel ntransistor 132 194 136 201 0 m9
rlabel ntransistor 132 183 136 190 0 m9
rlabel ntransistor 150 142 154 149 0 m7
rlabel ntransistor 132 166 136 173 0 m7
rlabel ntransistor 132 142 136 149 0 m8
rlabel ntransistor 150 166 154 173 0 m8
rlabel pwell 117 161 117 161 3 node4
rlabel pwell 117 154 117 154 3 node3
rlabel pwell 69 161 69 161 7 node5
rlabel pwell 69 154 69 154 7 node6
rlabel ntransistor 100 142 104 149 0 m6
rlabel ntransistor 82 166 86 173 0 m6
rlabel ntransistor 100 166 104 173 0 m5
rlabel ntransistor 82 142 86 149 0 m5
rlabel ntransistor 130 221 138 235 0 m12
rlabel ntransistor 101 221 105 235 0 m11
rlabel metal1 127 253 127 253 1 node15
rlabel ptransistor -19 267 173 269 0 m13
rlabel metal1 -11 86 -7 90 0 VDD
rlabel metal1 167 221 171 225 0 VSS
rlabel metal1 347 215 351 219 0 Vout
rlabel metal1 347 222 351 226 0 VSS
rlabel metal1 347 252 351 256 0 VDD
rlabel m2contact 29 134 29 134 1 node9
rlabel metal2 348 176 352 180 0 NBias
<< end >>
