magic
tech scmos
timestamp 695379491
<< polysilicon >>
rect -1 -27 4 27
<< metal1 >>
rect -2 23 5 28
<< labels >>
rlabel metal1 1 25 1 25 5 top
rlabel space 9 0 9 0 7 right
rlabel space -6 -1 -6 -1 3 left
rlabel polysilicon 1 -25 1 -25 1 bottom
<< end >>
